module dd1;
int random_number = $random;
inital begin ;
$display("Random number: %d", random_number);
end ;
endmodule; 